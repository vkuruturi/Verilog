module shifter_16bit (a, dir, shiftsize, out);
	input a;
	input dir;
	input shiftsize;

	output out;

	
endmodule
